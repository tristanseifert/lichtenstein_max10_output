LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY lichtenstein IS
      PORT(
			-- 24MHz main clock
			clkin:		  IN std_logic;
		
			-- SRAM bus
			sram_data: INOUT std_logic_vector(7 downto 0);
			sram_addr:   OUT std_logic_vector(17 downto 0);
			sram_oe:		 OUT std_logic;
			sram_ce:		 OUT std_logic;
			sram_we:		 OUT std_logic;
			
			-- SPI bus
			spi_cs:		  IN std_logic;
			spi_mosi:	  IN std_logic;
			spi_miso:	 OUT std_logic;
			spi_sck:		  IN std_logic;
			
			-- strobes from host
			ledout_en:	  IN std_logic;
			ledout_rst:	  IN std_logic;
			
			-- status outputs
			status:		 OUT std_logic_vector(2 downto 0);
			
			-- PWM output
			pwm_out:		 OUT std_logic_vector(15 downto 0)
		);
END lichtenstein;

ARCHITECTURE a OF lichtenstein IS

-- sram controller
component sram_controller
	PORT
	(
		-- clock and reset
		nreset:		IN STD_LOGIC;
		clk:			IN STD_LOGIC;
		
		-- SRAM bus
		address:		OUT STD_LOGIC_VECTOR(17 downto 0);
		data:			INOUT STD_LOGIC_VECTOR(7 downto 0);
		
		cs:			OUT STD_LOGIC := '1';
		oe:			OUT STD_LOGIC := '1';
		we:			OUT STD_LOGIC := '1';
		
		-- write interface
		wr_clk:		IN STD_LOGIC;
		wr_req:		IN STD_LOGIC := '1';
		wr_data:		IN STD_LOGIC_VECTOR(7 downto 0);
		wr_addr:		IN STD_LOGIC_VECTOR(17 downto 0);
		wr_full:		OUT STD_LOGIC;
		
		-- read interface
		rd_addr:		IN STD_LOGIC_VECTOR(17 downto 0);
		rd_data:		OUT STD_LOGIC_VECTOR(7 downto 0);
		rd_req:		IN STD_LOGIC := '0'
	);
end component;


-- SPI slave controller
component SPI_SLAVE is
    PORT (
        CLK      : in  std_logic; -- system clock
        RST      : in  std_logic; -- high active synchronous reset
        -- SPI SLAVE INTERFACE
        SCLK     : in  std_logic; -- SPI clock
        CS_N     : in  std_logic; -- SPI chip select, active in low
        MOSI     : in  std_logic; -- SPI serial data from master to slave
        MISO     : out std_logic; -- SPI serial data from slave to master
        -- USER INTERFACE
        DIN      : in  std_logic_vector(7 downto 0); -- input data for SPI master
        DIN_VLD  : in  std_logic; -- when DIN_VLD = 1, input data are valid
        READY    : out std_logic; -- when READY = 1, valid input data are accept
        DOUT     : out std_logic_vector(7 downto 0); -- output data from SPI master
        DOUT_VLD : out std_logic  -- when DOUT_VLD = 1, output data are valid
    );
end component;

-- command processor
component command_processor
	PORT
	(
		---------------------------------------
		-- clock and reset
		nreset:		IN STD_LOGIC;
		clk:			IN STD_LOGIC;
		
		---------------------------------------
		-- SPI interface
		spi_tx:		OUT STD_LOGIC_VECTOR(7 downto 0);
		spi_tx_valid:	OUT STD_LOGIC := '0';
		spi_tx_ready:	IN STD_LOGIC;
		
		spi_rx:		IN STD_LOGIC_VECTOR(7 downto 0);
		spi_rx_valid:	IN STD_LOGIC;
		
		---------------------------------------
		-- SRAM write interface
		sram_wr_data:	OUT STD_LOGIC_VECTOR(7 downto 0);
		sram_wr_addr:	OUT STD_LOGIC_VECTOR(17 downto 0);
		sram_wr_req:	OUT STD_LOGIC;
		sram_wr_full:	IN STD_LOGIC;
		
		---------------------------------------
		-- output registers
		out_addr:		OUT STD_LOGIC_VECTOR(17 downto 0);
		out_bytes:		OUT STD_LOGIC_VECTOR(15 downto 0);
		
		-- latch the addr/byte into one of the 16 output units
		out_latch:		OUT STD_LOGIC_VECTOR(15 downto 0)
	);
end component;

-- autogenerated component (mainpll.cmp)
component mainpll
	PORT
	(
		areset		: IN STD_LOGIC  := '0';
		inclk0		: IN STD_LOGIC  := '0';
		c0		: OUT STD_LOGIC ;
		c1		: OUT STD_LOGIC ;
		c2		: OUT STD_LOGIC ;
		locked		: OUT STD_LOGIC 
	);
end component;

-- output clocks from PLL
SIGNAL clk_24, clk_48, clk_800k	: std_logic;
SIGNAL pll_reset, pll_locked		: std_logic;

-- global reset, active 0
SIGNAL gReset							: std_logic := '1';

-- SRAM controller internal
signal sram_nreset					: std_logic;

-- SRAM write bus
signal sram_wrdata					: STD_LOGIC_VECTOR(7 downto 0);
signal sram_wraddr					: STD_LOGIC_VECTOR(17 downto 0);
signal sram_wrreq, sram_wrfull	: STD_LOGIC;

-- SRAM read bus
SIGNAL sram_rdaddr					: STD_LOGIC_VECTOR(17 downto 0);
SIGNAL sram_rddata					: STD_LOGIC_VECTOR(7 downto 0);
SIGNAL sram_rdreq						: STD_LOGIC := '0';

-- SPI interface
signal spi_reset						: STD_LOGIC := '0';

signal spi_tx							: STD_LOGIC_VECTOR(7 downto 0);
signal spi_tx_valid					: STD_LOGIC := '0';
signal spi_tx_ready					: STD_LOGIC;

signal spi_rx							: STD_LOGIC_VECTOR(7 downto 0);
signal spi_rx_valid					: STD_LOGIC;

-- command processor
signal cmd_nreset						: STD_LOGIC := '1';

-- output register bus
SIGNAL out_reg_addr					: STD_LOGIC_VECTOR(17 downto 0);
SIGNAL out_reg_bytes					: STD_LOGIC_VECTOR(15 downto 0);
SIGNAL out_reg_latch					: STD_LOGIC_VECTOR(15 downto 0);

BEGIN

-- instantiate main PLL
clocks: mainpll PORT MAP(areset => pll_reset, inclk0 => clkin, c0 => clk_24, 
	c1 => clk_48, c2 => clk_800k, locked => pll_locked
);

-- SRAM controller
sram: sram_controller PORT MAP(nreset => sram_nreset, clk => clk_48, 
	address => sram_addr, data => sram_data, cs => sram_ce, 
	oe => sram_oe, we => sram_we, wr_clk => clk_24, 
	wr_req => sram_wrreq, wr_data => sram_wrdata, 
	wr_addr => sram_wraddr, wr_full => sram_wrfull,
	rd_addr => sram_rdaddr, rd_data => sram_rddata, rd_req => sram_rdreq
);

-- SPI slave
spi: SPI_SLAVE PORT MAP(CLK => clk_48, RST => spi_reset, SCLK => spi_sck,
	CS_N => spi_cs, MOSI => spi_mosi, MISO => spi_miso, DIN => spi_tx,
	DIN_VLD => spi_tx_valid, READY => spi_tx_ready, DOUT => spi_rx,
	DOUT_VLD => spi_rx_valid
);

-- command processor
cmd: command_processor PORT MAP(nreset => cmd_nreset, clk => clk_48, 
	
	spi_tx => spi_tx, spi_tx_valid => spi_tx_valid, spi_rx => spi_rx,
	spi_tx_ready => spi_tx_ready,
	spi_rx_valid => spi_rx_valid, sram_wr_data => sram_wrdata, 
	
	sram_wr_addr => sram_wraddr, sram_wr_req => sram_wrreq,
	sram_wr_full => sram_wrfull,
	
	out_addr => out_reg_addr, out_bytes => out_reg_bytes, 
	out_latch => out_reg_latch
);



-- assert internal reset if external reset signal is asserted
PROCESS (clk_24) IS
BEGIN

	IF rising_edge(clk_24) THEN
		-- is the reset strobe asserted?
		IF ledout_rst = '0' THEN
			-- if so, assert reset
			gReset <= '0';
		ELSE
			-- de-assert reset
			gReset <= '1';
		END IF;
	END IF;
END PROCESS;

-- assert resets of all components if internal reset is asserted
PROCESS (clk_24) IS
BEGIN
	IF rising_edge(clk_24) THEN
		-- is reset low?
		IF gReset = '0' THEN
			-- if so, assert resets
			sram_nreset <= '0';
			cmd_nreset <= '0';

			spi_reset <= '1';
		ELSE
			-- de-assert resets
			sram_nreset <= '1';
			cmd_nreset <= '1';

			spi_reset <= '0';
		END IF;
	END IF;
END PROCESS;

END a;